* High Pass Filter Circuit
* Cutoff frequency: 1/(2*pi*R*C) = ~1.59kHz

* Input voltage source
V1 in 0 SIN(0 1 1k) AC 1

* High pass filter components
R1 in out 1k
C1 out 0 0.1uF

* Analysis commands
.tran 0.1ms 5ms
.print tran v(in) v(out)
.ac dec 10 10 100k
.print ac vdb(out) vp(out)
.end
